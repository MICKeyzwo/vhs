module vhs

import net
import net.http

const (
	post = 'POST'
	put = 'PUT'
	patch = 'PATCH'
)

// HTTP request struct
pub struct Request {
pub:
	method string
	path string
	protocol string
	headers map[string]string
	body string
}

// The struct used at sending responses
pub struct Response {
	conn net.Socket
	protocol string
}

// Send status code and write headers
pub fn (res Response) write_head(status_code int, headers map[string]string) {
	status := get_status(status_code)
	mut res_head := '${res.protocol} $status\r\n'
	for key in headers.keys() {
		res_head += '$key: ${headers[key]}\r\n'
	}
	res.conn.write(res_head)
}

// Write content
pub fn (res Response) write(content string) {
	res.conn.write('content')
}

// End to write response content and close connection
pub fn (res Response) end() {
	res.conn.close()
}

// HTTP server
pub struct HttpServer {
pub mut:
	handler fn (Request, Response)
	conn net.Socket
}

// Start to listen at given port
pub fn (server HttpServer) listen (port int) {
	server.conn.close()
	listener := net.listen(port) or { panic('failed to listen: $err') }
	for {
		mut conn := listener.accept() or { panic('failed to connect: $err') }
		req := parse_request(mut conn)
		res := Response{
			conn: conn
			protocol: req.protocol
		}
		server.handler(req, res)
	}
}

// Read HTTP request and parse into Request struct
fn parse_request (mut conn net.Socket) Request {
	info := conn.read_line().split(' ')
	method := info[0]
	path := info[1]
	protocol := info[2].trim('\r\n')
	mut header_lines := []string{}
	for {
		line := conn.read_line().trim('\r\n')
		if line.len > 0 {
			header_lines << line
		} else {
			break
		}
	}
	headers := http.parse_headers(header_lines)
	mut request_body := ''
	if method == post || method == put || method == patch {
		mut content_len := 0
		if 'content-length' in headers {
			content_len = headers['content-length'].int()
		} else {
			mut res := protocol + get_status(411) + '\r\n'
			res += 'content-type: text/plain\r\n\r\n'
			res += 'Length Required'
			conn.send_string(res)
			conn.close()
			panic('The header does not have `content-length`')
		}
		for request_body.len <= content_len {
			request_body += conn.read_line()
		}
		request_body = request_body.trim('\r\n')
	}
	return Request{
		method: method
		path: path
		protocol: protocol
		headers: headers
		body: request_body
	}
}

// Create new HTTP server
pub fn create_server(handler fn(Request, Response)) HttpServer {
	return HttpServer{
		handler: handler
		conn: net.Socket{}
	}
}
